`timescale 1ns/10ps

module  CONV(
            input		clk,
            input		reset,
            output	reg	busy,
            input		ready,

            output	reg [11:0]	iaddr,
            input	[19:0]	idata,

            output	reg 	cwr,
            output	reg [11:0] 	caddr_wr,
            output	reg [19:0] 	cdata_wr,

            output	reg 	crd,
            output	reg [11:0] 	caddr_rd,
            input	 [19:0]	cdata_rd,

            output	reg [2:0] 	csel
        );
reg [19:0] buffer[8:0];
reg [19:0] buffer_one[3:0];
reg [3:0] count;
reg [11:0] layerone_addr;
reg start = 1;
wire [19:0] com0, com1, max;
parameter k0 = 40'h000000a89e,
          k1 = 40'h00000092d5,
          k2 = 40'h0000006d43,
          k3 = 40'h0000001004,
          k4 = 40'hffffff8f71,
          k5 = 40'hffffff6e54,
          k6 = 40'hffffffa6d7,
          k7 = 40'hffffffc834,
          k8 = 40'hffffffac19;
wire [39:0] mul = {{20{buffer[0][19]}}, buffer[0]} * k0 + {{20{buffer[1][19]}}, buffer[1]} * k1 + {{20{buffer[2][19]}}, buffer[2]} * k2 + {{20{buffer[3][19]}}, buffer[3]} * k3 + {{20{buffer[4][19]}}, buffer[4]} * k4 + {{20{buffer[5][19]}}, buffer[5]} * k5 + {{20{buffer[6][19]}}, buffer[6]} * k6 + {{20{buffer[7][19]}}, buffer[7]} * k7 + {{20{buffer[8][19]}}, buffer[8]} * k8;
assign com0 = (buffer_one[0] >= buffer_one[1])?buffer_one[0]:buffer_one[1];
assign com1 = (buffer_one[2] >= buffer_one[3])?buffer_one[2]:buffer_one[3];
assign max = (com0 >= com1)?com0:com1;
integer i;
parameter bias = 20'h01310;

/*---------------------------------------------*/
always@(posedge clk or posedge reset) begin
    if(reset) begin
        busy <= 0;
        iaddr <= 1;
        cwr <= 0;
        caddr_wr <= 0;
        cdata_wr <= 0;
        crd <= 0;
        caddr_rd <= 0;
        csel <= 3'b001;
        count <= 0;
        buffer_one[0] <= 0;
        buffer_one[1] <= 0;
        buffer_one[2] <= 0;
        buffer_one[3] <= 0;
        layerone_addr <= 0;
        for(i = 0; i < 9; i = i + 1)
            buffer[i] <= 0;
    end
    else begin
        if(ready)
            busy <= 1;
        else begin
            if(start) begin
                start <= 0;
                busy <= 0;
            end
            else begin
                if(count == 12) begin
                    if(layerone_addr == 4030)
                        busy <= 0;
                    else
                        busy <= 1;
                end
                else
                    busy <= 1;
            end
        end
        case(count)
            /* layer 0 */
            0: begin
                if(ready)
                    iaddr <= iaddr;
                else begin
                    iaddr <= caddr_wr + 65;
                    buffer[5] <= idata;
                end
                count <= 1;
                if(caddr_wr[5:0] == 6'd0) begin //first col
                    buffer[0] <= 0;
                    buffer[3] <= 0;
                    buffer[6] <= 0;
                end
                else begin
                    buffer[0] <= buffer[1];
                    buffer[1] <= buffer[2];
                    buffer[3] <= buffer[4];
                    buffer[4] <= buffer[5];
                    buffer[6] <= buffer[7];
                    buffer[7] <= buffer[8];
                end
            end
            1: begin
                if(caddr_wr[5:0] == 6'd63) begin // final col
                    buffer[2] <= 0;
                    buffer[5] <= 0;
                    buffer[8] <= 0;
                    count <= 13;
                end
                else begin
                    if(caddr_wr >= 4032) begin
                        buffer[8] <= 0;
                    end
                    else begin
                        if(caddr_wr == 0) begin
                            buffer[5] <= idata;
                        end
                        else begin
                            buffer[8] <= idata;
                        end
                    end
                    if(caddr_wr <= 62) begin
                        if(caddr_wr == 0)
                            iaddr <= caddr_wr + 65;
                        else
                            iaddr <= caddr_wr;
                    end
                    else
                        iaddr <= caddr_wr - 63;
                    count <= 2;
                end
            end
            2: begin
                if(caddr_wr <= 62) begin //first row
                    if(caddr_wr == 0) begin
                        buffer[8] <= idata;
                        iaddr <= caddr_wr;
                        count <= 3;
                    end
                    else begin
                        count <= 13;
                    end
                end
                else begin //not first row
                    buffer[2] <= idata;
                    if(caddr_wr[5:0] == 6'd0) begin
                        count <= 4;
                        iaddr <= caddr_wr;
                    end
                    else
                        count <= 13;
                end
            end
            3: begin
                buffer[4] <= idata;
                iaddr <= caddr_wr + 64;
                count <= 4;
            end
            4: begin
                if(caddr_wr == 0) begin
                    buffer[7] <= idata;
                    count <= 13;
                end
                else begin
                    buffer[4] <= idata;
                    iaddr <= caddr_wr - 64;
                    count <= 5;
                end
            end
            5: begin
                buffer[1] <= idata;
                if(caddr_wr >= 4032) begin
                    buffer[7] <= 0;
                    count <= 13;
                end
                else begin
                    iaddr <= caddr_wr + 64;
                    count <= 6;
                end
            end
            6: begin
                buffer[7] <= idata;
                count <= 13;
            end
            /*  layer 1 */
            7: begin
                buffer_one[0] <= cdata_rd;
                caddr_rd <= layerone_addr + 1;
                count <= 8;
            end
            8: begin
                buffer_one[1] <= cdata_rd;
                caddr_rd <= layerone_addr + 64;
                count <= 9;
            end
            9: begin
                buffer_one[2] <= cdata_rd;
                caddr_rd <= layerone_addr + 65;
                count <= 10;
            end
            10: begin
                buffer_one[3] <= cdata_rd;
                caddr_rd <= layerone_addr + 2;
                count <= 11;
            end
            11: begin
                cwr <= 1;
                csel <= 3'b011;
                cdata_wr <= max;
                count <= 12;
            end
            12: begin
                cwr <= 0;
                csel <= 3'b001;
                caddr_wr <= caddr_wr + 1;
                if(layerone_addr[5:0] == 6'd62) begin
                    if(layerone_addr == 4030) begin
                        count <= 0;
                        caddr_wr <= 0;
                        iaddr <= 1;
                    end
                    else begin
                        layerone_addr <= layerone_addr + 66;
                        count <= 7;
                    end
                end
                else begin
                    layerone_addr <= layerone_addr + 2;
                    count <= 7;
                end
            end
            /* layer 0 output */
            13: begin
                cdata_wr <= mul[35:16] + mul[15] + bias;
                iaddr <= caddr_wr + 2;
                count <= 14;
            end
            14: begin
                cdata_wr <= (cdata_wr[19] == 1)?0:cdata_wr;
                cwr <= 1;
                count <= 15;
            end
            15: begin
                cwr <= 0;
                if(caddr_wr == 4095) begin
                    caddr_wr <= 0;
                    count <= 7;
                    crd <= 1;
                end
                else begin
                    caddr_wr <= caddr_wr + 1;
                    count <= 0;
                end
            end
        endcase
    end
end
endmodule
